
library IEEE;
use IEEE.STD_LOGIC_1164.all;

package prog_mem_content is

constant p_00 : std_logic_vector := X"1111";
constant p_01 : std_logic_vector := X"2222";
constant p_02 : std_logic_vector := X"3333";
constant p_03 : std_logic_vector := X"1234";
constant p_04 : std_logic_vector := X"1234";
constant p_05 : std_logic_vector := X"1234";
constant p_06 : std_logic_vector := X"1234";
constant p_07 : std_logic_vector := X"1234";
constant p_08 : std_logic_vector := X"1234";
constant p_09 : std_logic_vector := X"1234";
constant p_0A : std_logic_vector := X"1234";

end prog_mem_content;

